./bus/AdbBus.vhd